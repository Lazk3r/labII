library verilog;
use verilog.vl_types.all;
entity labII_vlg_vec_tst is
end labII_vlg_vec_tst;
