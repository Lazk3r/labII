lpm_counter4536_inst : lpm_counter4536 PORT MAP (
		aclr	 => aclr_sig,
		clk_en	 => clk_en_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
